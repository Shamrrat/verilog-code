module mux_condition(input i0,i1,s,output y);
assign y=s?i1:i0;
endmodule

