module top_module (
    input  clk,
    input  load,
    input  [511:0] data,
    output reg [511:0] q
);

    wire [511:0] left, right, next;

    // Neighbors with zero boundaries
    assign left  = {q[510:0], 1'b0};
    assign right = {1'b0, q[511:1]};

    // Rule 110 equation
    assign next = (q & ~right) | (left ^ q);

    always @(posedge clk) begin
        if (load)
            q <= data;
        else
            q <= next;
    end

endmodule
