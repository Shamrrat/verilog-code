module net_data;
wire a;
tri1 b;
wor  c;
wand d;
assign a=0;
assign a=1;
assign b=0;
assign c=0;
assign c=1;
assign d=0;
assign d=1;
initial
begin
 $display(" a=%b b=%b c=%b d=%b",a,b,c,d);
 end
endmodule
