 module default_value;
 wire a;
 wand b;
 wor c;
 supply1 d;
 supply0 e;
 tri0 f;
 tri1 g;
 reg i;
 integer j;
 time k;
 real l;
 realtime m;
 initial 
 begin 
 $display(" wire=%b wand=%b wor=%b supply1=%b supply0 =%b tri0=%b tri1=%b reg=%b integer=%d time=%t real=%f realtime=%f",a,b,c,d,e,f,g,i,j,k,l,m);
 end
 endmodule


