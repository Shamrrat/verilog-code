module memory;
reg [3:0] reg_a [0:2];
initial
begin
reg_a[0]=12;
reg_a[1]=10;
reg_a[2]=5;
$display("rega= %b  %d %h",reg_a[0],reg_a[1],reg_a[2]);
end
endmodule
