module and_gate(input wire a,b,output wire c);
and(c,a,b);
endmodule
