module top_module (
    input clk,
    input reset,
    input [31:0] in,
    output [31:0] out
);
        reg [31:0] in_d;  // previous-cycle input

    always @(posedge clk) begin
        if (reset) begin
            out  <= 32'b0;   // reset has priority
            in_d <= in;
        end else begin
            out  <= out | (in_d & ~in); // capture 1->0 transition
            in_d <= in;
        end
    end

endmodule
